module DramController_Verilog (
			input Clock,								// used to drive the state machine- stat changes occur on positive edge
			input Reset_L,     						// active low reset 
			input unsigned [12:0] Address,		// address bus from 68000
			input unsigned [15:0] DataIn,			// data bus in from 68000
			input DramSelect_L,     				// active low signal indicating dram is being addressed by 68000
			input WE_L,  								// active low write signal, otherwise assumed to be read
			input [1:0] BA ,

			output reg unsigned[15:0] DataOut, 				// data bus out to 68000
			output reg SDram_CKE_H,								// active high clock enable for dram chip
			output reg SDram_CS_L,								// active low chip select for dram chip
			output reg SDram_RAS_L,								// active low RAS select for dram chip
			output reg SDram_CAS_L,								// active low CAS select for dram chip		
			output reg SDram_WE_L,								// active low Write enable for dram chip
			output reg unsigned [12:0] SDram_Addr,			// 13 bit address bus dram chip	
			output reg unsigned [1:0] SDram_BA,				// 2 bit bank address
			input unsigned [15:0] 	SDram_DQ,			// 16 bit bi-directional data lines to dram chip
			
			output reg ResetOut_L,
			output reg LDQM,									
			output reg HDQM,
			output reg SDRAM_WE_L,								
	
			// Use only if you want to simulate dram controller state (e.g. for debugging)
			output reg [4:0] DramState
		); 	
		
		// WIRES and REGs
		
		reg  	[4:0] Command;										// 5 bit signal containing Dram_CKE_H, SDram_CS_L, SDram_RAS_L, SDram_CAS_L, SDram_WE_L
		reg [4:0] counter_re, counter_value;
		reg updateCounter, CounterLoad_H, CounterDone_H; 
		reg	TimerLoad_H ;										// logic 1 to load Timer on next clock
		reg   TimerDone_H ;										// set to logic 1 when timer reaches 0
		reg 	unsigned	[15:0] Timer;							// 16 bit timer value
		reg 	unsigned	[15:0] TimerValue;					// 16 bit timer preload value

		reg	RefreshTimerLoad_H;								// logic 1 to load refresh timer on next clock
		reg   RefreshTimerDone_H ;								// set to 1 when refresh timer reaches 0
		reg 	unsigned	[15:0] RefreshTimer;					// 16 bit refresh timer value
		reg 	unsigned	[15:0] RefreshTimerValue;			// 16 bit refresh timer preload value

		reg   unsigned [4:0] CurrentState;					// holds the current state of the dram controller
		reg   unsigned [4:0] NextState;						// holds the next state of the dram controller
		
		reg  	unsigned [1:0] BankAddress;
		reg  	unsigned [12:0] DramAddress;
		
		reg	DramDataLatch_H;									// used to indicate that data from SDRAM should be latched and held for 68000 after the CAS latency period
		reg  	unsigned [15:0]SDramWriteData;
		
		reg  FPGAWritingtoSDram_H;								// When '1' enables FPGA data out lines leading to SDRAM to allow writing, otherwise they are set to Tri-State "Z"
		reg  CPUReset_L;		
		reg  LDQM_O, HDQM_O;
		// 5 bit Commands to the SDRam

		parameter PoweringUp = 5'b00000 ;					// take CKE & CS low during power up phase, address and bank address = dont'care
		parameter DeviceDeselect  = 5'b11111;				// address and bank address = dont'care
		parameter NOP = 5'b10111;								// address and bank address = dont'care
		parameter BurstStop = 5'b10110;						// address and bank address = dont'care
		parameter ReadOnly = 5'b10101; 						// A10 should be logic 0, BA0, BA1 should be set to a value, other addreses = value
		parameter ReadAutoPrecharge = 5'b10101; 			// A10 should be logic 1, BA0, BA1 should be set to a value, other addreses = value
		parameter WriteOnly = 5'b10100; 						// A10 should be logic 0, BA0, BA1 should be set to a value, other addreses = value
		parameter WriteAutoPrecharge = 5'b10100 ;			// A10 should be logic 1, BA0, BA1 should be set to a value, other addreses = value
		parameter AutoRefresh = 5'b10001;
	
		parameter BankActivate = 5'b10011;					// BA0, BA1 should be set to a value, address A11-0 should be value
		parameter PrechargeSelectBank = 5'b10010;			// A10 should be logic 0, BA0, BA1 should be set to a value, other addreses = don't care
		
		parameter PrechargeAllBanks = 5'b10010;			// A10 should be logic 1, BA0, BA1 are dont'care, other addreses = don't care
		parameter ModeRegisterSet = 5'b10000;				// A10=0, BA1=0, BA0=0, Address = don't care
		parameter ExtModeRegisterSet = 5'b10000;			// A10=0, BA1=1, BA0=0, Address = value
		
	
		parameter InitialisingState = 5'h00;				// power on initialising state
		parameter WaitingForPowerUpState = 5'h01;		// waiting for power up state to complete
		parameter IssueFirstNOP = 5'h02;						// issuing 1st NOP after power up
		parameter PrechargingAllBanks = 5'h03;
		parameter Idle1 = 5'h04;
		parameter NOPAfterPrecharge = 5'h05;	
		parameter refresh_10 = 5'h06;
		parameter NOP_3x = 5'h07;
		parameter load_register = 5'h08;
		parameter waitNOP = 5'h09;
		parameter Issue3NOPS = 5'h0A;
		parameter Wait3NOP = 5'h0B;
		parameter SendRefresh = 5'h0C;		
		parameter PrechargeBanks = 5'h0D;
		parameter NOPAfterPrecharge_Re = 5'h0E;
		parameter IssueRefresh = 5'h0F;	
		parameter Issue3NOP    = 5'h10;
		parameter wait3NOP_Re = 5'h11;
		parameter IssueReadCommand = 5'h12;
		parameter waitUDS_LDS = 5'h13;
		parameter WaitCASLatency = 5'h14;
	        parameter Wait1Clock = 5'h15;
		parameter waitTerminate = 5'h16;		
		
		// TODO - Add your own states as per your own design
		

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// General Timer for timing and counting things: Loadable and counts down on each clock then produced a TimerDone signal and stops counting
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	always@(posedge Clock)
		if(TimerLoad_H == 1) 				// if we get the signal from another process to load the timer
			Timer <= TimerValue ;			// Preload timer
		else if(Timer != 16'd0) 			// otherwise, provided timer has not already counted down to 0, on the next rising edge of the clock		
			Timer <= Timer - 16'd1 ;		// subtract 1 from the timer value

	always@(Timer) begin
		TimerDone_H <= 0 ;					// default is not done
	
		if(Timer == 16'd0) 					// if timer has counted down to 0
			TimerDone_H <= 1 ;				// output '1' to indicate time has elapsed
	end

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Refresh Timer: Loadable and counts down on each clock then produces a RefreshTimerDone signal and stops counting
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

	always@(posedge Clock)
		if(RefreshTimerLoad_H == 1) 						// if we get the signal from another process to load the timer
			RefreshTimer  <= RefreshTimerValue ;		// Preload timer
		else if(RefreshTimer != 16'd0) 					// otherwise, provided timer has not already counted down to 0, on the next rising edge of the clock		
			RefreshTimer <= RefreshTimer - 16'd1 ;		// subtract 1 from the timer value

	always@(RefreshTimer) begin
		RefreshTimerDone_H <= 0 ;							// default is not done

		if(RefreshTimer == 16'd0) 								// if timer has counted down to 0
			RefreshTimerDone_H <= 1 ;						// output '1' to indicate time has elapsed
	end
	
	always@(posedge updateCounter)
		if(CounterLoad_H == 1) 				// if we get the signal from another process to load the timer
			counter_re <= counter_value ;			// Preload timer
		else if(counter_re != 16'd0) 			// otherwise, provided timer has not already counted down to 0, on the next rising edge of the clock		
			counter_re <= counter_re  - 16'd1 ;		// subtract 1 from the timer value

	always@(counter_re) begin
		CounterDone_H <= 0 ;					// default is not done
	
		if(counter_re == 16'd0) 					// if timer has counted down to 0
			CounterDone_H <= 1 ;				// output '1' to indicate time has elapsed
	end

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////-
// concurrent process state registers
// this process RECORDS the current state of the system.
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

   always@(posedge Clock, negedge Reset_L)
	begin
		if(Reset_L == 0) begin 							// asynchronous reset
			CurrentState <= InitialisingState ;
			ResetOut_L = 0;
		end	
		else 	begin									// state can change only on low-to-high transition of clock
			CurrentState <= NextState;		

			// these are the raw signals that come from the dram controller to the dram memory chip. 
			// This process expects the signals in the form of a 5 bit bus within the signal Command. The various Dram commands are defined above just beneath the architecture)

			SDram_CKE_H <= Command[4];			// produce the Dram clock enable
			SDram_CS_L  <= Command[3];			// produce the Dram Chip select
			SDram_RAS_L <= Command[2];			// produce the dram RAS
			SDram_CAS_L <= Command[1];			// produce the dram CAS
			SDram_WE_L  <= Command[0];			// produce the dram Write enable

			// Commands: 
			
			SDram_Addr <= DramAddress;		// output the row/column address to the dram
			SDram_BA   <= BankAddress;		// output the bank address to the dram

			// signals back to the 68000

			ResetOut_L 	<= CPUReset_L ;			// output the Reset out back to the 68000
			LDQM <=  LDQM_O;
			HDQM <=  HDQM_O;
			SDRAM_WE_L <= ~FPGAWritingtoSDram_H;
			
			// The signal FPGAWritingtoSDram_H can be driven by you when you need to turn on or tri-state the data bus out signals to the dram chip data lines DQ0-15
			// when you are reading from the dram you have to ensure they are tristated (so the dram chip can drive them)
			// when you are writing, you have to drive them to the value of SDramWriteData so that you 'present' your data to the dram chips
			// of course during a write, the dram WE signal will need to be driven low and it will respond by tri-stating its outputs lines so you can drive data in to it
			// remember the Dram chip has bi-directional data lines, when you read from it, it turns them on, when you write to it, it turns them off (tri-states them)

			if(FPGAWritingtoSDram_H == 1) 			// if CPU is doing a write, we need to turn on the FPGA data out lines to the SDRam and present Dram with CPU data 
			 SDram_DQ	<= SDramWriteData ;
			else
				SDram_DQ	<= 16'bZZZZZZZZZZZZZZZZ;
						// otherwise tri-state the FPGA data output lines to the SDRAM for anything other than writing to it
		
			DramState <= CurrentState ;					// output current state - useful for debugging so you can see you state machine changing states et
		end
	end	
	
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////-
// Concurrent process to Latch Data from Sdram after Cas Latency during read
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////-

// this process will latch whatever data is coming out of the dram data lines on the FALLING edge of the clock you have to drive DramDataLatch_H to logic 1
// remember there is a programmable CAS latency for the Zentel dram chip on the DE1 board it's 2 or 3 clock cycles which has to be programmed by you during the initialisation
// phase of the dram controller following a reset/power on
//
// During a read, after you have presented CAS command to the dram chip you will have to wait 2 clock cyles and then latch the data out here and present it back
// to the 68000 until the end of the 68000 bus cycles

	always@(negedge Clock)
	begin
		if(DramDataLatch_H == 1)      			// asserted during the read operation
			DataOut <= SDram_DQ ;					// store 16 bits of data regardless of width - don't worry about tri state since that will be handled by buffers outside dram controller
	end
	
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////-
// next state and output logic
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
	
	always@(*)
	begin
	
	// In Verilog/VHDL - you will recall - that combinational logic (i.e. logic with no storage) is created as long as you
	// provide a specific value for a signal in each and every possible path through a process
	// 
	// You can do this of course, but it gets tedious to specify a value for each signal inside every process state and every if-else test within those states
	// so the common way to do this is to define default values for all your signals and then override them with new values as and when you need to.
	// By doing this here, right at the start of a process, we ensure the compiler does not infer any storage for the signal, i.e. it creates
	// pure combinational logic (which is what we want)
	//
	// Let's start with default values for every signal and override as necessary, 
	//
	
		Command 	<= NOP ;												// assume no operation command for Dram chip
		NextState <= InitialisingState ;							// assume next state will always be idle state unless overridden the value used here is not important, we cimple have to assign something to prevent storage on the signal so anything will do
		
		TimerValue <= 16'h0000;										// no timer value 
		RefreshTimerValue <= 16'h0000 ;							// no refresh timer value
		TimerLoad_H <= 0;												// don't load Timer
		RefreshTimerLoad_H <= 0 ;									// don't load refresh timer
		DramAddress <= 13'h0000 ;									// no particular dram address
		BankAddress <= 2'b00 ;										// no particular dram bank address
		DramDataLatch_H <= 0;										// don't latch data yet
		SDramWriteData <= 16'h0000 ;								// nothing to write in particular
		CPUReset_L <= 0 ;												// default is reset to CPU (for the moment, though this will change when design is complete so that reset-out goes high at the end of the dram initialisation phase to allow CPU to resume)
		FPGAWritingtoSDram_H <= 0 ;								// default is to tri-state the FPGA data lines leading to bi-directional SDRam data lines, i.e. assume a read operation
		updateCounter  <= 1'b0;
		CounterLoad_H <= 0;
		counter_value <= 0;
		LDQM_O <=  1;
		HDQM_O <=  1;
		// put your current state/next state decision making logic here - here are a few states to get you started
		// during the initialising state, the drams have to power up and we cannot access them for a specified period of time (100 us)
		// we are going to load the timer above with a value equiv to 100us and then wait for timer to time out

// Begin initalization	
		if(CurrentState == InitialisingState ) begin
			TimerValue <= 16'h1338; // real value 1338									// chose a value equivalent to 100us at 50Mhz clock - you might want to shorten it to somthing small for simulation purposes
			TimerLoad_H <= 1 ;										// on next edge of clock, timer will be loaded and start to time out
			Command <= PoweringUp ;									// clock enable and chip select to the Zentel Dram chip must be held low (disabled) during a power up phase
			NextState <= WaitingForPowerUpState ;				// once we have loaded the timer, go to a new state where we wait for the 100us to elapse		
		end
		
		else if(CurrentState == WaitingForPowerUpState) begin
			Command <= PoweringUp ;									// no DRam clock enable or CS while witing for 100us timer
			
			if(TimerDone_H == 1) 									// if timer has timed out i.e. 100us have elapsed
				NextState <= IssueFirstNOP ;						// take CKE and CS to active and issue a 1st NOP command
			else
				NextState <= WaitingForPowerUpState ;			// otherwise stay here until power up time delay finished
		end
		
		else if(CurrentState == IssueFirstNOP) begin	 		// issue a valid NOP
			Command <= NOP ;											// send a valid NOP command to the dram chip
			NextState <= PrechargingAllBanks;
		end		
		
		else if(CurrentState ==  PrechargingAllBanks) begin
			Command <= PrechargeAllBanks;
			DramAddress <= 13'b00_10000000000;
			NextState <= NOPAfterPrecharge;
		end

		else if(CurrentState == NOPAfterPrecharge) begin
			counter_value <= 11;
			CounterLoad_H <= 1'b1;
			updateCounter <= 1'b1;
			Command <= NOP;
			DramAddress <= 13'h0;
			NextState <= refresh_10;
		end 
		else if (CurrentState == refresh_10) begin
		   updateCounter <= 1'b1;
		   if(CounterDone_H == 0) begin
			Command <= AutoRefresh;
			NextState <= NOP_3x;
		   end else if (CounterDone_H == 1) begin
		   	Command <= NOP;
			NextState <= load_register;
		   end
		end
		else if (CurrentState == NOP_3x) begin
			TimerValue <= 16'h0002;	
			TimerLoad_H <= 1;										
			Command <= NOP;									
			NextState <= waitNOP;
		end 
		else if (CurrentState == waitNOP) begin
			Command <= NOP;
			if(TimerDone_H == 1) begin 						
				NextState <= refresh_10 ;					
			end else
				NextState <= waitNOP ;			
		end
		else if (CurrentState == load_register) begin
			Command <= ModeRegisterSet;
			DramAddress <= 13'h220;
			NextState <= Issue3NOPS;
		end
		else if (CurrentState == Issue3NOPS) begin
			Command <= NOP;
			DramAddress <= 13'h0;
			NextState <= Wait3NOP;
			TimerValue <= 16'h0002;
			TimerLoad_H <= 1 ;
		end
		else if (CurrentState == Wait3NOP) begin
			Command <= NOP;
			if(TimerDone_H == 1) 									
				NextState <= SendRefresh ;						
			else
				NextState <= Wait3NOP ;
		end
		else if (CurrentState == SendRefresh) begin
			Command <= NOP;
			RefreshTimerLoad_H <= 1;
			RefreshTimerValue <= 16'h177; // 16'h177 is correct numer
			NextState <= Idle1;
		end
		// everything above above is just initalisation and setting the mode register to a value that is wanted: adjust CAS latency
		else if (CurrentState == Idle1) begin
			Command <= NOP;
			if(RefreshTimerDone_H)
			   NextState <= PrechargeBanks;
			else if ( (DramSelect_L == 0) && (AS_L == 0)) begin // this condition needs rto be changed. CHNAGE REQ
			    DramAddress <=  Address[12:0];
			    BankAddress <= BA[1:0]; // should bank address be part of address its self?
		            Command <= BankActivate; // activated the row  and the bank of DRAM
			    if (WE_L) 
				NextState <= IssueReadCommand; // if write enable_low is high then we should issue a read commmand
			   else 
				NextState <= waitUDS_LDS;
			end
			else
			NextState <= Idle1;
		end
// Handle the stupid refresh	
		else if (CurrentState == PrechargeBanks) begin
			Command <= PrechargeAllBanks;
			DramAddress <= 13'b000_10000000000;
			NextState <=  NOPAfterPrecharge_Re;
		end
		else if (CurrentState == NOPAfterPrecharge_Re) begin
			Command <= NOP;
			NextState <= IssueRefresh;
		end
		else if (CurrentState == IssueRefresh) begin 
			Command <= AutoRefresh;
			NextState <= Issue3NOP;
		end
		else if (CurrentState == Issue3NOP) begin
			TimerValue <= 16'h0002;	
			TimerLoad_H <= 1;										
			Command <= NOP;									
			NextState <= wait3NOP_Re;			
		end
		else if (CurrentState == wait3NOP_Re) begin
			Command <= NOP;
			if(TimerDone_H == 1) 									
				NextState <= SendRefresh ;						
			else
				NextState <= wait3NOP_Re ;	
		end
// BEGIN the stage of read and write states
		else if (CurrentState == IssueReadCommand) begin // CHANGE REQ: address selction
			DramAddress <= {3'b001, Address[9:0]};
			BankAddress <= BA[1:0];
			Command <= ReadAutoPrecharge;
			TimerValue <= 2;
			TimerLoad_H <= 1;
			NextState <= WaitCASLatency;
			LDQM_O <=  0;
			HDQM_O <=  0;
		end
		else if (CurrentState == WaitCASLatency) begin
			Command <= NOP;
			LDQM_O <=  0;
			HDQM_O <=  0;
			if(TimerDone_H) begin  
			  DramDataLatch_H <= 1; 
			  NextState <= waitTerminate;
			end 
			else 
			  NextState <= WaitCASLatency;
		end 
		else if (CurrentState == waitUDS_LDS) begin
			DramAddress <= {3'b001, Address[9:0]};
			BankAddress <= BA[1:0];
			LDQM_O <=  0;
			HDQM_O <=  0;
			Command <= WriteAutoPrecharge;
			FPGAWritingtoSDram_H <= 1;
			SDramWriteData <= DataIn;
			NextState <= Wait1Clock;
		end
		else if (CurrentState == Wait1Clock) begin
			Command <= NOP;
			LDQM_O <=  0;
			HDQM_O <=  0;
			FPGAWritingtoSDram_H <= 1;
			SDramWriteData <= DataIn;
			NextState <= waitTerminate;
		end
		else if (CurrentState == waitTerminate) begin
			Command <= NOP;
			NextState <= Idle1;
		end
		
	end	// always@ block
endmodule


